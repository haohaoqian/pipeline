`timescale 1ns / 1ps 
module InstructionMemory(Address, Instruction);
    input [31:0] Address;
    output reg [31:0] Instruction;

    always @(*)
    begin
        case ({1'b0,Address[30:2]})
            30'd0:  Instruction <= 32'h08000003;
            30'd1:  Instruction <= 32'h0800012f; 
            30'd2:  Instruction <= 32'h08000195; 
            30'd3:  Instruction <= 32'h0c000004; 
            30'd4:  Instruction <= 32'h3c017fff; 
            30'd5:  Instruction <= 32'h3428ffff; 
            30'd6:  Instruction <= 32'h03e8f824; 
            30'd7:  Instruction <= 32'h23ff001c; 
            30'd8:  Instruction <= 32'h3c014000; 
            30'd9:  Instruction <= 32'h34300000; 
            30'd10:  Instruction <= 32'h03e00008;
            30'd11:  Instruction <= 32'hae000008;
            30'd12:  Instruction <= 32'h3c01fffe;
            30'd13:  Instruction <= 32'h34287960;
            30'd14:  Instruction <= 32'hae080000;
            30'd15:  Instruction <= 32'hae080004;
            30'd16:  Instruction <= 32'h24040000;
            30'd17:  Instruction <= 32'h2408010a;
            30'd18:  Instruction <= 32'hac880000;
            30'd19:  Instruction <= 32'h24080342;
            30'd20:  Instruction <= 32'hac880004;
            30'd21:  Instruction <= 32'h240801a8;
            30'd22:  Instruction <= 32'hac880008;
            30'd23:  Instruction <= 32'h2408010b;
            30'd24:  Instruction <= 32'hac88000c;
            30'd25:  Instruction <= 32'h2408016c;
            30'd26:  Instruction <= 32'hac880010;
            30'd27:  Instruction <= 32'h2408009e;
            30'd28:  Instruction <= 32'hffffffff;
            30'd29:  Instruction <= 32'hac880014;
            30'd30:  Instruction <= 32'h2408017f;
            30'd31:  Instruction <= 32'hac880018;
            30'd32:  Instruction <= 32'h24080195;
            30'd33:  Instruction <= 32'hac88001c;
            30'd34:  Instruction <= 32'h24080269;
            30'd35:  Instruction <= 32'hac880020;
            30'd36:  Instruction <= 32'h240801d6;
            30'd37:  Instruction <= 32'hac880024;
            30'd38:  Instruction <= 32'h240803e5;
            30'd39:  Instruction <= 32'hac880028;
            30'd40:  Instruction <= 32'h240801ed;
            30'd41:  Instruction <= 32'hac88002c;
            30'd42:  Instruction <= 32'h240801ed;
            30'd43:  Instruction <= 32'hac880030;
            30'd44:  Instruction <= 32'h240801eb;
            30'd45:  Instruction <= 32'hac880034;
            30'd46:  Instruction <= 32'h2408037d;
            30'd47:  Instruction <= 32'hac880038;
            30'd48:  Instruction <= 32'h24080136;
            30'd49:  Instruction <= 32'hac88003c;
            30'd50:  Instruction <= 32'h24080023;
            30'd51:  Instruction <= 32'hac880040;
            30'd52:  Instruction <= 32'h24080324;
            30'd53:  Instruction <= 32'hac880044;
            30'd54:  Instruction <= 32'h24080095;
            30'd55:  Instruction <= 32'hac880048;
            30'd56:  Instruction <= 32'h240800ca;
            30'd57:  Instruction <= 32'hac88004c;
            30'd58:  Instruction <= 32'h24080361;
            30'd59:  Instruction <= 32'hac880050;
            30'd60:  Instruction <= 32'h240803dd;
            30'd61:  Instruction <= 32'hac880054;
            30'd62:  Instruction <= 32'h240800ba;
            30'd63:  Instruction <= 32'hac880058;
            30'd64:  Instruction <= 32'h2408014e;
            30'd65:  Instruction <= 32'hac88005c;
            30'd66:  Instruction <= 32'h240802f7;
            30'd67:  Instruction <= 32'hac880060;
            30'd68:  Instruction <= 32'h240801fb;
            30'd69:  Instruction <= 32'hac880064;
            30'd70:  Instruction <= 32'h24080032;
            30'd71:  Instruction <= 32'hac880068;
            30'd72:  Instruction <= 32'h240802cf;
            30'd73:  Instruction <= 32'hac88006c;
            30'd74:  Instruction <= 32'h240800a6;
            30'd75:  Instruction <= 32'hac880070;
            30'd76:  Instruction <= 32'h240802f9;
            30'd77:  Instruction <= 32'hac880074;
            30'd78:  Instruction <= 32'h240800e9;
            30'd79:  Instruction <= 32'hac880078;
            30'd80:  Instruction <= 32'h240803d7;
            30'd81:  Instruction <= 32'hac88007c;
            30'd82:  Instruction <= 32'h240801bd;
            30'd83:  Instruction <= 32'hac880080;
            30'd84:  Instruction <= 32'h24080007;
            30'd85:  Instruction <= 32'hac880084;
            30'd86:  Instruction <= 32'h24080061;
            30'd87:  Instruction <= 32'hac880088;
            30'd88:  Instruction <= 32'h24080005;
            30'd89:  Instruction <= 32'hac88008c;
            30'd90:  Instruction <= 32'h240802aa;
            30'd91:  Instruction <= 32'hac880090;
            30'd92:  Instruction <= 32'h2408035d;
            30'd93:  Instruction <= 32'hac880094;
            30'd94:  Instruction <= 32'h24080166;
            30'd95:  Instruction <= 32'hac880098;
            30'd96:  Instruction <= 32'h240802df;
            30'd97:  Instruction <= 32'hac88009c;
            30'd98:  Instruction <= 32'h24080336;
            30'd99:  Instruction <= 32'hac8800a0;
            30'd100:  Instruction <= 32'h2408021e;
            30'd101:  Instruction <= 32'hac8800a4;
            30'd102:  Instruction <= 32'h240801c7;
            30'd103:  Instruction <= 32'hac8800a8;
            30'd104:  Instruction <= 32'h24080392;
            30'd105:  Instruction <= 32'hac8800ac;
            30'd106:  Instruction <= 32'h2408011d;
            30'd107:  Instruction <= 32'hac8800b0;
            30'd108:  Instruction <= 32'h240803d0;
            30'd109:  Instruction <= 32'hac8800b4;
            30'd110:  Instruction <= 32'h24080058;
            30'd111:  Instruction <= 32'hac8800b8;
            30'd112:  Instruction <= 32'h2408031b;
            30'd113:  Instruction <= 32'hac8800bc;
            30'd114:  Instruction <= 32'h24080065;
            30'd115:  Instruction <= 32'hac8800c0;
            30'd116:  Instruction <= 32'h240803af;
            30'd117:  Instruction <= 32'hac8800c4;
            30'd118:  Instruction <= 32'h240801b1;
            30'd119:  Instruction <= 32'hac8800c8;
            30'd120:  Instruction <= 32'h240803b0;
            30'd121:  Instruction <= 32'hac8800cc;
            30'd122:  Instruction <= 32'h24080109;
            30'd123:  Instruction <= 32'hac8800d0;
            30'd124:  Instruction <= 32'h240801d2;
            30'd125:  Instruction <= 32'hac8800d4;
            30'd126:  Instruction <= 32'h240800e7;
            30'd127:  Instruction <= 32'hac8800d8;
            30'd128:  Instruction <= 32'h240803d8;
            30'd129:  Instruction <= 32'hac8800dc;
            30'd130:  Instruction <= 32'h2408036d;
            30'd131:  Instruction <= 32'hac8800e0;
            30'd132:  Instruction <= 32'h24080308;
            30'd133:  Instruction <= 32'hac8800e4;
            30'd134:  Instruction <= 32'h24080217;
            30'd135:  Instruction <= 32'hac8800e8;
            30'd136:  Instruction <= 32'h24080366;
            30'd137:  Instruction <= 32'hac8800ec;
            30'd138:  Instruction <= 32'h240802b3;
            30'd139:  Instruction <= 32'hac8800f0;
            30'd140:  Instruction <= 32'h24080003;
            30'd141:  Instruction <= 32'hac8800f4;
            30'd142:  Instruction <= 32'h24080180;
            30'd143:  Instruction <= 32'hac8800f8;
            30'd144:  Instruction <= 32'h24080168;
            30'd145:  Instruction <= 32'hac8800fc;
            30'd146:  Instruction <= 32'h24080156;
            30'd147:  Instruction <= 32'hac880100;
            30'd148:  Instruction <= 32'h240800f3;
            30'd149:  Instruction <= 32'hac880104;
            30'd150:  Instruction <= 32'h240801d9;
            30'd151:  Instruction <= 32'hac880108;
            30'd152:  Instruction <= 32'h240802c6;
            30'd153:  Instruction <= 32'hac88010c;
            30'd154:  Instruction <= 32'h2408003e;
            30'd155:  Instruction <= 32'hac880110;
            30'd156:  Instruction <= 32'h24080222;
            30'd157:  Instruction <= 32'hac880114;
            30'd158:  Instruction <= 32'h240801d2;
            30'd159:  Instruction <= 32'hac880118;
            30'd160:  Instruction <= 32'h24080330;
            30'd161:  Instruction <= 32'hac88011c;
            30'd162:  Instruction <= 32'h240802ee;
            30'd163:  Instruction <= 32'hac880120;
            30'd164:  Instruction <= 32'h24080046;
            30'd165:  Instruction <= 32'hac880124;
            30'd166:  Instruction <= 32'h24080261;
            30'd167:  Instruction <= 32'hac880128;
            30'd168:  Instruction <= 32'h24080243;
            30'd169:  Instruction <= 32'hac88012c;
            30'd170:  Instruction <= 32'h240801b5;
            30'd171:  Instruction <= 32'hac880130;
            30'd172:  Instruction <= 32'h24080171;
            30'd173:  Instruction <= 32'hac880134;
            30'd174:  Instruction <= 32'h2408013d;
            30'd175:  Instruction <= 32'hac880138;
            30'd176:  Instruction <= 32'h240801a8;
            30'd177:  Instruction <= 32'hac88013c;
            30'd178:  Instruction <= 32'h240802f8;
            30'd179:  Instruction <= 32'hac880140;
            30'd180:  Instruction <= 32'h2408033f;
            30'd181:  Instruction <= 32'hac880144;
            30'd182:  Instruction <= 32'h2408032b;
            30'd183:  Instruction <= 32'hac880148;
            30'd184:  Instruction <= 32'h24080351;
            30'd185:  Instruction <= 32'hac88014c;
            30'd186:  Instruction <= 32'h24080037;
            30'd187:  Instruction <= 32'hac880150;
            30'd188:  Instruction <= 32'h24080105;
            30'd189:  Instruction <= 32'hac880154;
            30'd190:  Instruction <= 32'h2408023a;
            30'd191:  Instruction <= 32'hac880158;
            30'd192:  Instruction <= 32'h2408033d;
            30'd193:  Instruction <= 32'hac88015c;
            30'd194:  Instruction <= 32'h2408030d;
            30'd195:  Instruction <= 32'hac880160;
            30'd196:  Instruction <= 32'h2408034a;
            30'd197:  Instruction <= 32'hac880164;
            30'd198:  Instruction <= 32'h240802b8;
            30'd199:  Instruction <= 32'hac880168;
            30'd200:  Instruction <= 32'h240801ba;
            30'd201:  Instruction <= 32'hac88016c;
            30'd202:  Instruction <= 32'h24080228;
            30'd203:  Instruction <= 32'hac880170;
            30'd204:  Instruction <= 32'h240802c6;
            30'd205:  Instruction <= 32'hac880174;
            30'd206:  Instruction <= 32'h240800c5;
            30'd207:  Instruction <= 32'hac880178;
            30'd208:  Instruction <= 32'h240800f1;
            30'd209:  Instruction <= 32'hac88017c;
            30'd210:  Instruction <= 32'h2408034e;
            30'd211:  Instruction <= 32'hac880180;
            30'd212:  Instruction <= 32'h24080313;
            30'd213:  Instruction <= 32'hac880184;
            30'd214:  Instruction <= 32'h240803bb;
            30'd215:  Instruction <= 32'hac880188;
            30'd216:  Instruction <= 32'h240800f6;
            30'd217:  Instruction <= 32'hac88018c;
            30'd218:  Instruction <= 32'h24080267;
            30'd219:  Instruction <= 32'hac880190;
            30'd220:  Instruction <= 32'h24080083;
            30'd221:  Instruction <= 32'hac880194;
            30'd222:  Instruction <= 32'h240801a8;
            30'd223:  Instruction <= 32'hac880198;
            30'd224:  Instruction <= 32'h2408001c;
            30'd225:  Instruction <= 32'hac88019c;
            30'd226:  Instruction <= 32'h2408004e;
            30'd227:  Instruction <= 32'hac8801a0;
            30'd228:  Instruction <= 32'h24080165;
            30'd229:  Instruction <= 32'hac8801a4;
            30'd230:  Instruction <= 32'h24080019;
            30'd231:  Instruction <= 32'hac8801a8;
            30'd232:  Instruction <= 32'h240800e4;
            30'd233:  Instruction <= 32'hac8801ac;
            30'd234:  Instruction <= 32'h2408006c;
            30'd235:  Instruction <= 32'hac8801b0;
            30'd236:  Instruction <= 32'h2408038e;
            30'd237:  Instruction <= 32'hac8801b4;
            30'd238:  Instruction <= 32'h24080389;
            30'd239:  Instruction <= 32'hac8801b8;
            30'd240:  Instruction <= 32'h2408011f;
            30'd241:  Instruction <= 32'hac8801bc;
            30'd242:  Instruction <= 32'h240802df;
            30'd243:  Instruction <= 32'hac8801c0;
            30'd244:  Instruction <= 32'h24080340;
            30'd245:  Instruction <= 32'hac8801c4;
            30'd246:  Instruction <= 32'h24080314;
            30'd247:  Instruction <= 32'hac8801c8;
            30'd248:  Instruction <= 32'h24080184;
            30'd249:  Instruction <= 32'hac8801cc;
            30'd250:  Instruction <= 32'h2408025c;
            30'd251:  Instruction <= 32'hac8801d0;
            30'd252:  Instruction <= 32'h240803d5;
            30'd253:  Instruction <= 32'hac8801d4;
            30'd254:  Instruction <= 32'h240801a0;
            30'd255:  Instruction <= 32'hac8801d8;
            30'd256:  Instruction <= 32'h240803e1;
            30'd257:  Instruction <= 32'hac8801dc;
            30'd258:  Instruction <= 32'h240800f0;
            30'd259:  Instruction <= 32'hac8801e0;
            30'd260:  Instruction <= 32'h240801e2;
            30'd261:  Instruction <= 32'hac8801e4;
            30'd262:  Instruction <= 32'h240801de;
            30'd263:  Instruction <= 32'hac8801e8;
            30'd264:  Instruction <= 32'h2408039b;
            30'd265:  Instruction <= 32'hac8801ec;
            30'd266:  Instruction <= 32'h24080240;
            30'd267:  Instruction <= 32'hac8801f0;
            30'd268:  Instruction <= 32'h24080018;
            30'd269:  Instruction <= 32'hac8801f4;
            30'd270:  Instruction <= 32'h24080051;
            30'd271:  Instruction <= 32'hac8801f8;
            30'd272:  Instruction <= 32'h24080008;
            30'd273:  Instruction <= 32'hac8801fc;
            30'd274:  Instruction <= 32'h8e160014;
            30'd275:  Instruction <= 32'h24110080;
            30'd276:  Instruction <= 32'h24120000;
            30'd277:  Instruction <= 32'h24130000;
            30'd278:  Instruction <= 32'h0251502a;
            30'd279:  Instruction <= 32'h1140000e;
            30'd280:  Instruction <= 32'h2253ffff;
            30'd281:  Instruction <= 32'h0660000a;
            30'd282:  Instruction <= 32'h00135080;
            30'd283:  Instruction <= 32'h008a5020;
            30'd284:  Instruction <= 32'h8d4b0000;
            30'd285:  Instruction <= 32'h8d4c0004;
            30'd286:  Instruction <= 32'h018b682a;
            30'd287:  Instruction <= 32'h11a00004;
            30'd288:  Instruction <= 32'had4c0000;
            30'd289:  Instruction <= 32'had4b0004;
            30'd290:  Instruction <= 32'h2273ffff;
            30'd291:  Instruction <= 32'h08000119;
            30'd292:  Instruction <= 32'h22520001;
            30'd293:  Instruction <= 32'h08000116;
            30'd294:  Instruction <= 32'h8e170014;
            30'd295:  Instruction <= 32'h240800ff;
            30'd296:  Instruction <= 32'hae08000c;
            30'd297:  Instruction <= 32'h02f6b822;
            30'd298:  Instruction <= 32'h24080003;
            30'd299:  Instruction <= 32'hae080008;
            30'd300:  Instruction <= 32'h24150000;
            30'd301:  Instruction <= 32'h24160000;
            30'd302:  Instruction <= 32'h0800012e;
            30'd303:  Instruction <= 32'h24080001;
            30'd304:  Instruction <= 32'hae080008;
            30'd305:  Instruction <= 32'h12a00006;
            30'd306:  Instruction <= 32'h24010001;
            30'd307:  Instruction <= 32'h12a10007;
            30'd308:  Instruction <= 32'h24010002;
            30'd309:  Instruction <= 32'h12a10009;
            30'd310:  Instruction <= 32'h24010003;
            30'd311:  Instruction <= 32'h12a1000b;
            30'd312:  Instruction <= 32'h24140100;
            30'd313:  Instruction <= 32'h32e9000f;
            30'd314:  Instruction <= 32'h08000146;
            30'd315:  Instruction <= 32'h24140200;
            30'd316:  Instruction <= 32'h32e900f0;
            30'd317:  Instruction <= 32'h00094902;
            30'd318:  Instruction <= 32'h08000146;
            30'd319:  Instruction <= 32'h24140400;
            30'd320:  Instruction <= 32'h32e90f00;
            30'd321:  Instruction <= 32'h00094a02;
            30'd322:  Instruction <= 32'h08000146;
            30'd323:  Instruction <= 32'h24140800;
            30'd324:  Instruction <= 32'h32e9f000;
            30'd325:  Instruction <= 32'h00094b02;
            30'd326:  Instruction <= 32'h24010000;
            30'd327:  Instruction <= 32'h1121001e;
            30'd328:  Instruction <= 32'h24010001;
            30'd329:  Instruction <= 32'h1121001e;
            30'd330:  Instruction <= 32'h24010002;
            30'd331:  Instruction <= 32'h1121001e;
            30'd332:  Instruction <= 32'h24010003;
            30'd333:  Instruction <= 32'h1121001e;
            30'd334:  Instruction <= 32'h24010004;
            30'd335:  Instruction <= 32'h1121001e;
            30'd336:  Instruction <= 32'h24010005;
            30'd337:  Instruction <= 32'h1121001e;
            30'd338:  Instruction <= 32'h24010006;
            30'd339:  Instruction <= 32'h1121001e;
            30'd340:  Instruction <= 32'h24010007;
            30'd341:  Instruction <= 32'h1121001e;
            30'd342:  Instruction <= 32'h24010008;
            30'd343:  Instruction <= 32'h1121001e;
            30'd344:  Instruction <= 32'h24010009;
            30'd345:  Instruction <= 32'h1121001e;
            30'd346:  Instruction <= 32'h2401000a;
            30'd347:  Instruction <= 32'h1121001e;
            30'd348:  Instruction <= 32'h2401000b;
            30'd349:  Instruction <= 32'h1121001e;
            30'd350:  Instruction <= 32'h2401000c;
            30'd351:  Instruction <= 32'h1121001e;
            30'd352:  Instruction <= 32'h2401000d;
            30'd353:  Instruction <= 32'h1121001e;
            30'd354:  Instruction <= 32'h2401000e;
            30'd355:  Instruction <= 32'h1121001e;
            30'd356:  Instruction <= 32'h2401000f;
            30'd357:  Instruction <= 32'h1121001e;
            30'd358:  Instruction <= 32'h369400c0;
            30'd359:  Instruction <= 32'h08000185;
            30'd360:  Instruction <= 32'h369400f9;
            30'd361:  Instruction <= 32'h08000185;
            30'd362:  Instruction <= 32'h369400a4;
            30'd363:  Instruction <= 32'h08000185;
            30'd364:  Instruction <= 32'h369400b0;
            30'd365:  Instruction <= 32'h08000185;
            30'd366:  Instruction <= 32'h36940099;
            30'd367:  Instruction <= 32'h08000185;
            30'd368:  Instruction <= 32'h36940092;
            30'd369:  Instruction <= 32'h08000185;
            30'd370:  Instruction <= 32'h36940082;
            30'd371:  Instruction <= 32'h08000185;
            30'd372:  Instruction <= 32'h369400f8;
            30'd373:  Instruction <= 32'h08000185;
            30'd374:  Instruction <= 32'h36940080;
            30'd375:  Instruction <= 32'h08000185;
            30'd376:  Instruction <= 32'h36940090;
            30'd377:  Instruction <= 32'h08000185;
            30'd378:  Instruction <= 32'h36940088;
            30'd379:  Instruction <= 32'h08000185;
            30'd380:  Instruction <= 32'h36940083;
            30'd381:  Instruction <= 32'h08000185;
            30'd382:  Instruction <= 32'h369400c6;
            30'd383:  Instruction <= 32'h08000185;
            30'd384:  Instruction <= 32'h369400a1;
            30'd385:  Instruction <= 32'h08000185;
            30'd386:  Instruction <= 32'h36940086;
            30'd387:  Instruction <= 32'h08000185;
            30'd388:  Instruction <= 32'h3694008e;
            30'd389:  Instruction <= 32'h24010004;
            30'd390:  Instruction <= 32'h22b50001;
            30'd391:  Instruction <= 32'hae140010;
            30'd392:  Instruction <= 32'h16a10009;
            30'd393:  Instruction <= 32'h22d60001;
            30'd394:  Instruction <= 32'h24010005;
            30'd395:  Instruction <= 32'h24150000;
            30'd396:  Instruction <= 32'h16c10005;
            30'd397:  Instruction <= 32'hae000008;
            30'd398:  Instruction <= 32'hae00000c;
            30'd399:  Instruction <= 32'h24080fff;
            30'd400:  Instruction <= 32'hae080010;
            30'd401:  Instruction <= 32'h03400008;
            30'd402:  Instruction <= 32'h24080003;
            30'd403:  Instruction <= 32'hae080008;
            30'd404:  Instruction <= 32'h03400008;
            30'd405:  Instruction <= 32'h00000000;
            30'd406:  Instruction <= 32'h00000000;
            30'd407:  Instruction <= 32'h00000000;
            30'd408:  Instruction <= 32'h03400008;
            default:  Instruction <= 32'h00000000;
        endcase
    end

endmodule